module angleFP2Int(
	input [15:0] angle,
	output [15:0] int
	);