module HalfPrecesion2Int(
	input [15:0] angleFP,
	output [15:0] angleInt
	);
	
	always@(*) begin
	
	end
endmodule 