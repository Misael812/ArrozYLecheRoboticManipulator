module tb_angleFP2CyclesPositive;

endmodule 